
----------------------------------------------------
--defining our packages
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package GLOBAL is
	constant data_bus_width: 		integer := 16;
	constant addr_bus_width: 		integer := 8;
	constant control_bus_width: 	integer := 6;
	constant register_adr_width: 	integer := 4;
	constant register_addr_width: integer := 4;	
	type register_block is array (0 to (register_addr_width - 1) ) of std_logic_vector( (data_bus_width - 1) downto 0 );
	type ram_type is array (0 to (addr_bus_width - 1) ) of std_logic_vector( (data_bus_width - 1) downto 0 );
end GLOBAL;

-----------------------------------------------------

--ALU 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
entity alu is
 Port ( inp_a : in signed(7 downto 0);
 inp_b : in signed(7 downto 0);
 sel : in STD_LOGIC_VECTOR (2 downto 0);
 out_alu : out signed(7 downto 0));
end alu;

architecture Behavioral of alu is
begin
process(inp_a, inp_b, sel) 
begin
case sel is
 when "000" => 
 out_alu<= inp_a + inp_b; 
 when "001" => 
 out_alu<= inp_a - inp_b;
 when "010" => 
 out_alu<= inp_a - 1; 
 when "011" => 
 out_alu<= inp_a + 1; 
 when "100" => 
 out_alu<= inp_a and inp_b;
 when "101" => 
 out_alu<= inp_a or inp_b;
 when "110" => 
 out_alu<= not inp_a ;
 when "111" => 
 out_alu<= inp_a xor inp_b;
 when others =>
 NULL;
end case;
 
end process; 

end Behavioral;

-------------------------------------
--Data path 
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use WORK.GLOBAL.ALL;

entity data_path is
	port	(	
				CS: 			in 	std_logic;
				OPERAND:		in		std_logic_vector( (register_addr_width - 1) downto 0 );
				DIN: 			in 	std_logic_vector( (addr_bus_width - 1) downto 0 );	
				DOUT: 		out 	std_logic_vector( (data_bus_width - 1) downto 0 );
				CLK:			in		std_logic;
				INSTRUCTION:in		std_logic_vector( 1 downto 0)
			);
end data_path;


Architecture implement of data_path is
		signal latched_operand: std_logic_vector( (data_bus_width - 1) downto 0 ) := (others => '0');
		signal registers : register_block;
		--signal inp_b_sliced : std_logic_vector(7 downto 0);
		--signal control : std_logic_vector(2 downto 0); 


--component alu is
--  port (
 --   inp_a   : in std_logic_vector(7 downto 0);
 --   inp_b   : in std_logic_vector(7 downto 0);
   -- sel     : in std_logic_vector(2 downto 0);
  --  out_alu : out std_logic_vector(7 downto 0)
 -- );
--end component alu;
	
begin
--control <= '0' &  INSTRUCTION;
data_alu: process( CLK , CS , OPERAND , INSTRUCTION , DIN ) is

  begin
    if rising_edge( CLK ) AND CS = '1' then
      case INSTRUCTION is
			when "00" =>
			   -- latch OPERAND
				latched_operand <= registers( conv_integer( OPERAND ) ); 
			when "01" =>
			   --add latched operand to OPERAND
				latched_operand <= latched_operand + registers( conv_integer( OPERAND ) );
			when "10" =>
				--put OPERAND on DOUT
				DOUT <= registers( conv_integer( OPERAND ) );
			when "11" =>
				--set OPERAND to DIN
				registers( conv_integer( OPERAND ))(15 downto 8)  <= DIN;
			when others =>
      end case;
    end if;
 end process data_alu;
--inp_b_sliced <= registers(conv_integer(OPERAND))(15 downto 8); 

--  alu_inst : alu
 --   port map (
  --    inp_a   => std_logic_vector(latched_operand(7 downto 0)),
   --   inp_b   => inp_b_sliced,
    --  sel     => control,
     -- out_alu => DOUT(7 downto 0)
    --);

end implement;

------------------------------------
--counter
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use WORK.GLOBAL.ALL;

entity counter is port 
		(
			CLK: 	in 	std_logic;
			CS:	in		std_logic;
			DOUT:	out 	std_logic_vector( (addr_bus_width - 1) downto 0 )
		); 
end counter;

architecture counter_core of counter is
	signal counter_variable: std_logic_vector( (addr_bus_width - 1) downto 0 ) := (others => '0');
begin

	counting: process ( CLK , CS )
	begin
		if rising_edge( CLK ) AND CS = '1' then
			DOUT <= counter_variable;
			counter_variable <= counter_variable + 1;
		end if;
	end process;
end counter_core;

----------------------------------------------
--Conttrol unit
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use WORK.GLOBAL.ALL;

entity control_unit is port 
		(
			CLOCK: 			in 	std_logic;
			DATA_BUS: 		inout std_logic_vector( (data_bus_width - 1) downto 0 );
			CONTROL_BUS:	inout std_logic_vector( (control_bus_width - 1) downto 0 );
			IR: 				inout std_logic_vector( (control_bus_width - 1) downto 0 );
			MAR: 				inout std_logic_vector( (addr_bus_width - 1) downto 0 );
			MDR: 				inout	std_logic_vector( (data_bus_width - 1) downto 0 )
		); 
end control_unit;

architecture control_core of control_unit is
	
	component counter is port 
	(
		CLK: 	in 	std_logic;
		CS:	in		std_logic;
		DOUT:	out 	std_logic_vector( (addr_bus_width - 1) downto 0 )
	);
	end component;
		
	component data_path is port	
	(	
		CS: 			in 	std_logic;
		OPERAND:		in		std_logic_vector( (register_addr_width - 1) downto 0 );
		DIN: 			in 	std_logic_vector( (addr_bus_width - 1) downto 0 );	
		DOUT: 		out 	std_logic_vector( (data_bus_width - 1) downto 0 );
		CLK:			in		std_logic;
		INSTRUCTION:in		std_logic_vector( 1 downto 0)
	);
	end component;
	
	begin
	
	program_counter: counter port map 
	(
		CLK => CLOCK,
		CS => CONTROL_BUS(0),
		DOUT => MAR
	);

	alu: data_path port map
	(
		CLK => CLOCK,
		INSTRUCTION => CONTROL_BUS(2 downto 1), 
		OPERAND => CONTROL_BUS(5 downto 2),
		CS =>  CONTROL_BUS(5),
		DIN => MAR,
		DOUT => MDR
	);

end control_core;
--------------------------------------------------------------------
---memory block 

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.Numeric_Std.all;
use WORK.GLOBAL.ALL;

entity memory_block is
	port	(	
				ADDR: in 	std_logic_vector( (addr_bus_width - 1) downto 0 );
				DIN:	in		std_logic_vector( (data_bus_width - 1) downto 0 );
				DOUT: out 	std_logic_vector( (data_bus_width - 1) downto 0 );	
				CLK:	in		std_logic;
				RW:	in		std_logic; -- 0 = read, 1 = write
				CS0:	in 	std_logic;
				CS1:	in 	std_logic
			);
end memory_block;

Architecture cell of memory_block is
	signal ram : ram_type;
begin

memory_process: process( CLK , DIN , ADDR , RW , CS0 , CS1) is
  begin
    if rising_edge( CLK ) AND CS0 = '1' AND CS1 = '1' then
		case RW is
			when '0' => --read 
				DOUT <= ram( conv_integer( ADDR ) );
			when '1' => --write 
				ram( conv_integer( ADDR ) ) <= DIN;
				DOUT <= "ZZZZZZZZZZZZZZZZ"; -- TODO: tri-state is hardcoded, should be generic	
			when others =>
				DOUT <= "ZZZZZZZZZZZZZZZZ"; -- TODO: tri-state is hardcoded, should be generic
		end case;
    end if;
 end process memory_process;
end cell;

----------------------------------------------------------------------------------------------
---Alu testbench 
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
  
ENTITY Tb_alu IS
END Tb_alu;
  
ARCHITECTURE behavior OF Tb_alu IS
   
 COMPONENT alu
 PORT(
 inp_a : IN signed(7 downto 0);
 inp_b : IN signed(7 downto 0);
 sel : IN std_logic_vector(2 downto 0);
 out_alu : OUT signed(7 downto 0)
 );
 END COMPONENT;
  
 signal inp_a : signed(7 downto 0) := (others => '0');
 signal inp_b : signed(7 downto 0) := (others => '0');
 signal sel : std_logic_vector(2 downto 0) := (others => '0');
 signal out_alu : signed(7 downto 0);
 
BEGIN
 uut: alu PORT MAP (
 inp_a => inp_a,
 inp_b => inp_b,
 sel => sel,
 out_alu => out_alu
 );
 

 stim_proc: process
 begin

 wait for 100 ns;

 inp_a <= "00001001";
 inp_b <= "00001111";
 sel <= "111";
 end process;
END;
----------------------------------------------------------------------------------------
--MAIN CODE 
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use WORK.GLOBAL.ALL;

entity main is port 
		(
			CLOCK: in std_logic
		); 
end main;

architecture computer of main is
	signal memory_request: std_logic;
	signal read_write: std_logic;
	signal addr_bus: std_logic_vector( (addr_bus_width - 1) downto 0 );
	signal data_bus: std_logic_vector( (data_bus_width - 1) downto 0 );
	signal control_bus: std_logic_vector( (control_bus_width - 1) downto 0 );	
	signal instruction_register: std_logic_vector( (control_bus_width - 1) downto 0 );
	signal memory_address_register: std_logic_vector( (addr_bus_width - 1) downto 0 );
	signal memory_data_register: std_logic_vector( (data_bus_width - 1) downto 0 );
	
	component memory_block port 
	(
		ADDR: in 	std_logic_vector( (addr_bus_width - 1) downto 0 );
		DIN:	in		std_logic_vector( (data_bus_width - 1) downto 0 );
		DOUT: out 	std_logic_vector( (data_bus_width - 1) downto 0 );	
		CLK:	in		std_logic;
		RW:	in		std_logic; 
		CS0:	in 	std_logic;
		CS1:	in 	std_logic
	);
	end component;
	
	component control_unit port 
	(
		CLOCK: 			in 	std_logic;
		DATA_BUS: 		in 	std_logic_vector( (data_bus_width - 1) downto 0 );
		CONTROL_BUS:	out 	std_logic_vector( (control_bus_width - 1) downto 0 );
		IR: 				inout std_logic_vector( (control_bus_width - 1) downto 0 );
		MAR: 				inout std_logic_vector( (addr_bus_width - 1) downto 0 );
		MDR: 				inout	std_logic_vector( (data_bus_width - 1) downto 0 )
	); 
	end component;
	signal mycs1 :std_logic; 
	begin
	mycs1 <= not addr_bus(3);
	M1: memory_block port map 
	(
		ADDR => addr_bus,
		DIN => data_bus,
		DOUT => data_bus,
		CLK => CLOCK,
		RW => read_write,
		CS0 => memory_request,
		CS1 => mycs1
	);

	M2: memory_block port map
	(
		ADDR => addr_bus,
		DIN => data_bus,
		DOUT =>  data_bus,
		CLK => CLOCK,
		RW => read_write,
		CS0 => memory_request,
		CS1 => addr_bus(3)
	);
	
	CU: control_unit port map 
	(
		CLOCK => CLOCK,
		DATA_BUS => data_bus,
		CONTROL_BUS => control_bus,
		IR => instruction_register,
		MAR => memory_address_register,
		MDR => memory_data_register
	);
	
end computer;


----------------
---main code testbench 
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use WORK.GLOBAL.ALL;

entity main_tb is
end main_tb;

architecture tb_architecture of main_tb is
    constant addr_bus_width: integer := 8; -- Update with appropriate width
    constant data_bus_width: integer := 8; -- Update with appropriate width
    constant control_bus_width: integer := 8; -- Update with appropriate width

    signal CLOCK: std_logic := '0';
    signal memory_request: std_logic;
    signal read_write: std_logic;
    signal addr_bus: std_logic_vector((addr_bus_width - 1) downto 0);
    signal data_bus: std_logic_vector((data_bus_width - 1) downto 0);
    signal control_bus: std_logic_vector((control_bus_width - 1) downto 0);
    signal instruction_register: std_logic_vector((control_bus_width - 1) downto 0);
    signal memory_address_register: std_logic_vector((addr_bus_width - 1) downto 0);
    signal memory_data_register: std_logic_vector((data_bus_width - 1) downto 0);

    component main
        port (
            CLOCK: in std_logic
        );
    end component;

    component memory_block
        port (
            ADDR: in std_logic_vector((addr_bus_width - 1) downto 0);
            DIN: in std_logic_vector((data_bus_width - 1) downto 0);
            DOUT: out std_logic_vector((data_bus_width - 1) downto 0);
            CLK: in std_logic;
            RW: in std_logic;
            CS0: in std_logic;
            CS1: in std_logic
        );
    end component;

    component control_unit
        port (
            CLOCK: in std_logic;
            DATA_BUS: in std_logic_vector((data_bus_width - 1) downto 0);
            CONTROL_BUS: out std_logic_vector((control_bus_width - 1) downto 0);
            IR: inout std_logic_vector((control_bus_width - 1) downto 0);
            MAR: inout std_logic_vector((addr_bus_width - 1) downto 0);
            MDR: inout std_logic_vector((data_bus_width - 1) downto 0)
        );
    end component;

    signal mycs1 :std_logic; 

begin

    UUT: main port map (CLOCK => CLOCK);

    mycs1 <= not addr_bus(3);
    
    M1: memory_block port map 
    (
        ADDR => addr_bus,
        DIN => data_bus,
        DOUT => data_bus,
        CLK => CLOCK,
        RW => read_write,
        CS0 => memory_request,
        CS1 => mycs1
    );

    M2: memory_block port map
    (
        ADDR => addr_bus,
        DIN => data_bus,
        DOUT => data_bus,
        CLK => CLOCK,
        RW => read_write,
        CS0 => memory_request,
        CS1 => addr_bus(3)
    );
    
    CU: control_unit port map 
    (
        CLOCK => CLOCK,
        DATA_BUS => data_bus,
        CONTROL_BUS => control_bus,
        IR => instruction_register,
        MAR => memory_address_register,
        MDR => memory_data_register
    );

    -- Clock process
    process
    begin
        while now < 100 ns loop -- Update simulation time if necessary
            CLOCK <= '0';
            wait for 5 ns; -- Update clock period if necessary
            CLOCK <= '1';
            wait for 5 ns; -- Update clock period if necessary
        end loop;
        wait;
    end process;

end tb_architecture;

-----------------------

--cpu FSM approach : 



library ieee;
use ieee.std_logic_1164.all ;
use ieee. std_logic_unsigned.all ;

entity CPU8BIT2 is
port ( data: inout std_logic_vector (7 downto 0);
adress: out std_logic_vector(5 downto 0);
oe: out std_logic;
we: out std_logic ;
rst : in std_logic;
clk : in std_logic);

end;
 architecture CPU_ARCH of CPU8BIT2 is
signal akku: std_logic_vector(8 downto 0); 
signal adreg:  std_logic_vector(5 downto 0);
signal pc: std_logic_vector (5 downto 0);
signal states : std_logic_vector(2 downto 0);
begin
process(clk,rst)
begin
if ( rst = '0') then
adreg <= (others => '0'); 
states <= "000";
akku <= (others => '0');
pc <= (others => '0');
elsif rising_edge (clk) then

if ( states = "000") then
pc <= adreg + 1;
adreg <= data(5 downto 0);
else
 adreg <= pc;
end if;

case states is

when "010" => akku <= ("0" & akku(7 downto 0)) + ("0" & data); 
when "011" => akku(7 downto 0) <= akku(7 downto 0) nor data; 
when "101" => akku(8) <= '0'; 
when others => null; --instr. fetch, jcc taken (000), sta (001)
end case;

--State machine
if ( states /= "000") then states <= "000"; 
elsif (data(7 downto 6) = "11" and akku(8)='1') then states <= "101";
else states <= "0" & not data(7 downto 6); 
 end if;
end if;
end process;

adress <= adreg;
data <= "ZZZZZZZZ" when states /= "001" else akku(7 downto 0);
oe <= '1' when (clk='1' or states = "001" or rst='0' or states = "101") else '0';
we <= '1' when (clk='1' or states /= "001" or rst='0') else '0';
end CPU_ARCH;

--testbench 
library ieee;
use ieee.std_logic_1164.all;

entity CPU8BIT2_Test is
end entity;

architecture tb_arch of CPU8BIT2_Test is
    component CPU8BIT2 is
        port (
            data   : inout std_logic_vector(7 downto 0);
            adress : out std_logic_vector(5 downto 0);
            oe     : out std_logic;
            we     : out std_logic;
            rst    : in std_logic;
            clk    : in std_logic
        );
    end component;

    signal data_tb   : std_logic_vector(7 downto 0) := (others => '0');
    signal adress_tb : std_logic_vector(5 downto 0) := (others => '0');
    signal oe_tb     : std_logic := '0';
    signal we_tb     : std_logic := '0';
    signal rst_tb    : std_logic := '0';
    signal clk_tb    : std_logic := '0';

begin

    uut: CPU8BIT2
    port map(
        data   => data_tb,
        adress => adress_tb,
        oe     => oe_tb,
        we     => we_tb,
        rst    => rst_tb,
        clk    => clk_tb
    );

clk_process: process
  begin
    while now < 10000 ns loop
      clk_tb <= '0';
      wait for 10 ns;
      clk_tb <= '1';
      wait for 10 ns;
    end loop;
    wait;
  end process;

    stimulus_proc: process
    begin
        -- Initialize inputs
        rst_tb <= '1';
         wait for 10 ns; 
	data_tb <= "00000000" ;
	wait for 10 ns; 
	data_tb <= "01000100" ;
	wait for 10 ns; 
	data_tb <= "10100000";
        wait; -- Wait indefinitely
    end process;

    -- Add assertions or checks if required

end architecture;
